`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: sustech
// Engineer: happys
// 
// Create Date: 2020/12/09 11:16:04
// Design Name: SnakeGame
// Module Name: snake
// Project Name: VGA
//////////////////////////////////////////////////////////////////////////////////


module snake();
endmodule
